module Mem (
    input clk, 
    input MemRead, 
    input MemWrite, 
    input [7:0] addr, 
    input [31:0] data_in, 
    input [2:0]func3, 
    output reg [31:0] data_out
    );
 reg [7:0] mem [0:255];
 //assign data_out = {mem[addr+3], mem[addr+2],mem[addr+1],mem[addr] };

  always @(posedge clk) begin
 data_out <= {mem[addr+3], mem[addr+2],mem[addr+1],mem[addr] };
 end

 always@ (negedge clk) begin
  if (MemRead)begin
  if (func3==3'b000) data_out<={{24{mem[addr][7]}},mem[addr]};//lb
  if (func3==3'b001) data_out<={{16{mem[addr+1][7]}},mem[addr+1], mem[addr]};//lh
  if (func3==3'b010) data_out<={mem[addr+3], mem[addr+2],mem[addr+1],mem[addr] };//lw
  if (func3==3'b100) data_out<={{24{1'b0}},mem[addr]};//lbu
  if (func3==3'b101) data_out<={{16{1'b0}},mem[addr+1], mem[addr]};//lhu
  end
   if(MemWrite)begin
 if (func3==3'b000) mem[addr]<=data_in[7:0];
 if (func3==3'b001) {mem[addr+1], mem[addr]}<=data_in[15:0];
 if (func3==3'b010) {mem[addr+3], mem[addr+2],mem[addr+1],mem[addr] }<=data_in;
 end
 end
 initial begin/*
mem[0]=32'h00002283;// lw x5, 0(x0)
mem[1]=32'h00402b03;// lw x22, 4(x0)
mem[2]=32'h00802b83;// lw x23, 8(x0)
mem[3]=32'h41628333;// sub x6, x5, x22
mem[4]=32'h0042e093;// ori x1, x5, 4
mem[5]=32'h002b1513;// Loop: slli x10, x22, 2
mem[6]=32'h01950533;// add x10, x10, x25
mem[7]=32'h00032483;//lw x9, 0(x6)
mem[8]=32'h000063b7;// lui x7, 6
mem[9]=32'h00004417;// auipc x8, 4
mem[10]=32'h030003e7;// jalr x7, 48(x0)
mem[11]=32'h04001a63;// bne x0, x0, Exit
mem[12]=32'h001b0b13;// addi x22, x22, 1
mem[13]=32'h035a8663;// beq x21, x21, label
mem[14]=32'h00c0036f;// jal x6, branch
mem[15]=32'h022c8263;// beq x25, x2, label
mem[16]=32'h02219063;// bne x3, x2, label
mem[17]=32'h001b4e63;// branch: blt x22, x1, label
mem[18]=32'h0021dc63;// bge x3, x2, label
mem[19]=32'h0021ea63;// bltu x3, x2, label
mem[20]=32'h0021f863;// bgeu x3, x2, label
mem[21]=32'h00528503;// lb x10, 5(x5)
mem[22]=32'h00529503;// lh x10, 5(x5)
mem[23]=32'h0052a503;// lw x10, 5(x5)
mem[24]=32'h0043c503;// label: lbu x10, 4(x7)
mem[25]=32'h0092d503;// lhu x10, 9(x5)
mem[26]=32'h00110523;// sb x1, 10(x2)
mem[27]=32'h00a10183;// lb x3, 10(x2)
mem[28]=32'h00711523;// sh x7, 10(x2)
mem[29]=32'h00410093;// addi x1, x2, 4
mem[30]=32'h00412093;// slti x1, x2, 4
mem[31]=32'h00413093;// sltiu x1, x2, 4
mem[32]=32'h00458503;// Exit: lb x10, 4(x11)
mem[33]=32'h003100b3;// add x1, x2, x3
mem[34]=32'h403100b3;//sub x1, x2, x3
mem[35]=32'h003110b3;// sll x1, x2, x3
mem[36]=32'h003120b3;// slt x1, x2, x3
mem[37]=32'h00712523;// sw x7, 10(x2)
mem[38]=32'h00414093;// xori x1, x2, 4
mem[38]=32'h00416093;// ori x1, x2, 4
mem[39]=32'h00417093;// andi x1, x2, 4
mem[40]=32'h002c9293;// slli x5, x25, 2
mem[41]=32'h002cd293;// srli x5, x25, 2
mem[42]=32'h4022dc93;// srai x25, x5, 2
mem[43]=32'h003130b3;// sltu x1, x2, x3
mem[44]=32'h003140b3;// xor x1, x2, x3
mem[45]=32'h003150b3;// srl x1, x2, x3
mem[46]=32'h403150b3;// sra x1, x2, x3
mem[47]=32'h003160b3;// or x1, x2, x3
mem[48]=32'h003170b3;// and x1, x2, x3
mem[49]=32'h00100073;//  ebreak
mem[50]=32'h00000033;// add x0, x0, x0
mem[51]=32'h40938333 ;//sub x6, x7, x9
mem[52]=32'h0110000f;//  fence 1, 1
mem[53]=32'h00000073;// ecall*/
//{mem[3],mem[2],mem[1],mem[0]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 //added to be skipped since PC starts with 4 after reset
 {mem[3],mem[2],mem[1],mem[0]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[7],mem[6],mem[5],mem[4]}=32'h0c802083;//32'b000000000000_00000_010_00001_0000011 ; //lw x1, 0(x0)
 {mem[11],mem[10],mem[9],mem[8]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[15],mem[14],mem[13],mem[12]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[19],mem[18],mem[17],mem[16]} = 32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[23],mem[22],mem[21],mem[20]} = 32'h0cc02103;//32'b000000000100_00000_010_00010_0000011 ; //lw x2, 4(x0)
 {mem[27],mem[26],mem[25],mem[24]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[31],mem[30],mem[29],mem[28]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[35],mem[34],mem[33],mem[32]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[39],mem[38],mem[37],mem[36]}=32'h0d002183;//32'b000000001000_00000_010_00011_0000011 ; //lw x3, 8(x0)
 {mem[43],mem[42],mem[41],mem[40]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[47],mem[46],mem[45],mem[44]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[51],mem[50],mem[49],mem[48]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[55],mem[54],mem[53],mem[52]}=32'b0000000_00010_00001_110_00100_0110011 ; //or x4, x1, x2
 {mem[59],mem[58],mem[57],mem[56]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[63],mem[62],mem[61],mem[60]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[67],mem[66],mem[65],mem[64]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[71],mem[70],mem[69],mem[68]}=32'b0_000001_00011_00100_000_0000_0_1100011; //beq x4, x3, 16
 {mem[75],mem[74],mem[73],mem[72]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[79],mem[78],mem[77],mem[76]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[83],mem[82],mem[81],mem[80]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[87],mem[86],mem[85],mem[84]}=32'b0000000_00010_00001_000_00011_0110011 ; //add x3, x1, x2
 {mem[91],mem[90],mem[89],mem[88]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[95],mem[94],mem[93],mem[92]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[99],mem[98],mem[97],mem[96]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[103],mem[102],mem[101],mem[100]}=32'b0000000_00010_00011_000_00101_0110011 ; //add x5, x3, x2
 {mem[107],mem[106],mem[105],mem[104]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[111],mem[110],mem[109],mem[108]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0 
 {mem[115],mem[114],mem[113],mem[112]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[119],mem[118],mem[117],mem[116]}=32'h0c502a23;//32'b0000000_00101_00000_010_01100_0100011; //sw x5, 12(x0)
 {mem[123],mem[122],mem[121],mem[120]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[127],mem[126],mem[125],mem[124]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[131],mem[130],mem[129],mem[128]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[135],mem[134],mem[133],mem[132]}=32'b000000001100_00000_010_00110_0000011 ; //lw x6, 12(x0)
 {mem[139],mem[138],mem[137],mem[136]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[143],mem[142],mem[141],mem[140]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[147],mem[146],mem[145],mem[144]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[151],mem[150],mem[149],mem[148]}=32'b0000000_00001_00110_111_00111_0110011 ; //and x7, x6, x1
 {mem[155],mem[154],mem[153],mem[152]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[159],mem[158],mem[157],mem[156]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[163],mem[162],mem[161],mem[160]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[167],mem[166],mem[165],mem[164]}=32'b0100000_00010_00001_000_01000_0110011 ; //sub x8, x1, x2
 {mem[171],mem[170],mem[169],mem[168]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[175],mem[174],mem[173],mem[172]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[179],mem[178],mem[177],mem[176]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[183],mem[182],mem[181],mem[180]}=32'b0000000_00010_00001_000_00000_0110011 ; //add x0, x1, x2
 {mem[187],mem[186],mem[185],mem[184]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[191],mem[190],mem[189],mem[188]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[195],mem[194],mem[193],mem[192]}=32'b0000000_00000_00000_000_00000_0110011 ; //add x0, x0, x0
 {mem[199],mem[198],mem[197],mem[196]}=32'b0000000_00001_00000_000_01001_0110011 ; //add x9, x0, x1
  mem[200]=8'd17;
  mem[201]=8'd0; 
  mem[202]=8'd0; 
  mem[203]=8'd0; 
  mem[204]=8'd9; 
  mem[205]=8'd0; 
  mem[206]=8'd0;
  mem[207]=8'd0; 
  mem[208]=8'd25; 
  mem[209]=8'd0;
  mem[210]=8'd0;
  mem[211]=8'd0;
  mem[212]=8'd25;
  mem[213]=8'd0;  
  mem[214]=8'd0;  
  mem[215]=8'b00000001;  
  mem[216]=8'b01100000; //24577 for 15-16
  mem[217]=8'b10101010;//170, -86
 end 
endmodule